// Broderick Bownds & Sebastian Heredia
// brbownds@g.hmc.edu & dheredia@g.hmc.edu
// November 18, 2025

// twiddle_vectors.sv contains the LUT for twiddle vectors used for a 512-point FFT.

module twiddle_vectors
  #(parameter bit_width = 16, N = 512, M = 9)
  
  (input logic clk, reset,
   input logic [M - 1:0] twiddle_adr,
   output logic [2*bit_width - 1:0] twiddle_out);
  
  logic [2*bit_width - 1:0] twiddle [0:(N/2) - 1];      // "256 twiddles of size 32-bits each"
    
  // Indexing k from 0 to 255 for a 512-point FFT:
    assign twiddle[0]   = 32'h7FFF0000; // cos: 1.000000, sin:0.000000
    assign twiddle[1]   = 32'h7FFD0192; // cos: 0.999925, sin:0.012272
    assign twiddle[2]   = 32'h7FF50324; // cos: 0.999699, sin:0.024541
    assign twiddle[3]   = 32'h7FE904B6; // cos: 0.999322, sin:0.036807
    assign twiddle[4]   = 32'h7FD80648; // cos: 0.998795, sin:0.049068
    assign twiddle[5]   = 32'h7FC107D9; // cos: 0.998118, sin:0.061321
    assign twiddle[6]   = 32'h7FA6096A; // cos: 0.997290, sin:0.073565
    assign twiddle[7]   = 32'h7F860AFB; // cos: 0.996313, sin:0.085797
    assign twiddle[8]   = 32'h7F610C8C; // cos: 0.995185, sin:0.098017
    assign twiddle[9]   = 32'h7F370E1C; // cos: 0.993907, sin:0.110222
    assign twiddle[10]  = 32'h7F090FAB; // cos: 0.992480, sin:0.122411
    assign twiddle[11]  = 32'h7ED5113A; // cos: 0.990903, sin:0.134581
    assign twiddle[12]  = 32'h7E9C12C8; // cos: 0.989177, sin:0.146730
    assign twiddle[13]  = 32'h7E5F1455; // cos: 0.987301, sin:0.158858
    assign twiddle[14]  = 32'h7E1D15E2; // cos: 0.985278, sin:0.170962
    assign twiddle[15]  = 32'h7DD5176E; // cos: 0.983105, sin:0.183040
    assign twiddle[16]  = 32'h7D8918F9; // cos: 0.980785, sin:0.195090
    assign twiddle[17]  = 32'h7D391A82; // cos: 0.978317, sin:0.207111
    assign twiddle[18]  = 32'h7CE31C0B; // cos: 0.975702, sin:0.219101
    assign twiddle[19]  = 32'h7C881D93; // cos: 0.972940, sin:0.231058
    assign twiddle[20]  = 32'h7C291F1A; // cos: 0.970031, sin:0.242980
    assign twiddle[21]  = 32'h7BC5209F; // cos: 0.966976, sin:0.254866
    assign twiddle[22]  = 32'h7B5C2223; // cos: 0.963776, sin:0.266713
    assign twiddle[23]  = 32'h7AEE23A6; // cos: 0.960431, sin:0.278520
    assign twiddle[24]  = 32'h7A7C2528; // cos: 0.956940, sin:0.290285
    assign twiddle[25]  = 32'h7A0526A8; // cos: 0.953306, sin:0.302006
    assign twiddle[26]  = 32'h79892826; // cos: 0.949528, sin:0.313682
    assign twiddle[27]  = 32'h790929A3; // cos: 0.945607, sin:0.325310
    assign twiddle[28]  = 32'h78842B1F; // cos: 0.941544, sin:0.336890
    assign twiddle[29]  = 32'h77FA2C99; // cos: 0.937339, sin:0.348419
    assign twiddle[30]  = 32'h776B2E11; // cos: 0.932993, sin:0.359895
    assign twiddle[31]  = 32'h76D82F87; // cos: 0.928506, sin:0.371317
    assign twiddle[32]  = 32'h764130FB; // cos: 0.923880, sin:0.382683
    assign twiddle[33]  = 32'h75A5326E; // cos: 0.919114, sin:0.393992
    assign twiddle[34]  = 32'h750433DF; // cos: 0.914210, sin:0.405241
    assign twiddle[35]  = 32'h745F354D; // cos: 0.909168, sin:0.416430
    assign twiddle[36]  = 32'h73B536BA; // cos: 0.903989, sin:0.427555
    assign twiddle[37]  = 32'h73073824; // cos: 0.898674, sin:0.438616
    assign twiddle[38]  = 32'h7254398C; // cos: 0.893224, sin:0.449611
    assign twiddle[39]  = 32'h719D3AF2; // cos: 0.887640, sin:0.460539
    assign twiddle[40]  = 32'h70E23C56; // cos: 0.881921, sin:0.471397
    assign twiddle[41]  = 32'h70223DB8; // cos: 0.876070, sin:0.482184
    assign twiddle[42]  = 32'h6F5E3F17; // cos: 0.870087, sin:0.492898
    assign twiddle[43]  = 32'h6E964073; // cos: 0.863973, sin:0.503538
    assign twiddle[44]  = 32'h6DC941CE; // cos: 0.857729, sin:0.514103
    assign twiddle[45]  = 32'h6CF84325; // cos: 0.851355, sin:0.524590
    assign twiddle[46]  = 32'h6C23447A; // cos: 0.844854, sin:0.534998
    assign twiddle[47]  = 32'h6B4A45CD; // cos: 0.838225, sin:0.545325
    assign twiddle[48]  = 32'h6A6D471C; // cos: 0.831470, sin:0.555570
    assign twiddle[49]  = 32'h698B4869; // cos: 0.824589, sin:0.565732
    assign twiddle[50]  = 32'h68A649B4; // cos: 0.817585, sin:0.575808
    assign twiddle[51]  = 32'h67BC4AFB; // cos: 0.810457, sin:0.585798
    assign twiddle[52]  = 32'h66CF4C3F; // cos: 0.803208, sin:0.595699
    assign twiddle[53]  = 32'h65DD4D81; // cos: 0.795837, sin:0.605511
    assign twiddle[54]  = 32'h64E84EBF; // cos: 0.788346, sin:0.615232
    assign twiddle[55]  = 32'h63EE4FFB; // cos: 0.780737, sin:0.624859
    assign twiddle[56]  = 32'h62F15133; // cos: 0.773010, sin:0.634393
    assign twiddle[57]  = 32'h61F05268; // cos: 0.765167, sin:0.643832
    assign twiddle[58]  = 32'h60EB539B; // cos: 0.757209, sin:0.653173
    assign twiddle[59]  = 32'h5FE354C9; // cos: 0.749136, sin:0.662416
    assign twiddle[60]  = 32'h5ED755F5; // cos: 0.740951, sin:0.671559
    assign twiddle[61]  = 32'h5DC7571D; // cos: 0.732654, sin:0.680601
    assign twiddle[62]  = 32'h5CB35842; // cos: 0.724247, sin:0.689541
    assign twiddle[63]  = 32'h5B9C5964; // cos: 0.715731, sin:0.698376
    assign twiddle[64]  = 32'h5A825A82; // cos: 0.707107, sin:0.707107
    assign twiddle[65]  = 32'h59645B9C; // cos: 0.698376, sin:0.715731
    assign twiddle[66]  = 32'h58425CB3; // cos: 0.689541, sin:0.724247
    assign twiddle[67]  = 32'h571D5DC7; // cos: 0.680601, sin:0.732654
    assign twiddle[68]  = 32'h55F55ED7; // cos: 0.671559, sin:0.740951
    assign twiddle[69]  = 32'h54C95FE3; // cos: 0.662416, sin:0.749136
    assign twiddle[70]  = 32'h539B60EB; // cos: 0.653173, sin:0.757209
    assign twiddle[71]  = 32'h526861F0; // cos: 0.643832, sin:0.765167
    assign twiddle[72]  = 32'h513362F1; // cos: 0.634393, sin:0.773010
    assign twiddle[73]  = 32'h4FFB63EE; // cos: 0.624859, sin:0.780737
    assign twiddle[74]  = 32'h4EBF64E8; // cos: 0.615232, sin:0.788346
    assign twiddle[75]  = 32'h4D8165DD; // cos: 0.605511, sin:0.795837
    assign twiddle[76]  = 32'h4C3F66CF; // cos: 0.595699, sin:0.803208
    assign twiddle[77]  = 32'h4AFB67BC; // cos: 0.585798, sin:0.810457
    assign twiddle[78]  = 32'h49B468A6; // cos: 0.575808, sin:0.817585
    assign twiddle[79]  = 32'h4869698B; // cos: 0.565732, sin:0.824589
    assign twiddle[80]  = 32'h471C6A6D; // cos: 0.555570, sin:0.831470
    assign twiddle[81]  = 32'h45CD6B4A; // cos: 0.545325, sin:0.838225
    assign twiddle[82]  = 32'h447A6C23; // cos: 0.534998, sin:0.844854
    assign twiddle[83]  = 32'h43256CF8; // cos: 0.524590, sin:0.851355
    assign twiddle[84]  = 32'h41CE6DC9; // cos: 0.514103, sin:0.857729
    assign twiddle[85]  = 32'h40736E96; // cos: 0.503538, sin:0.863973
    assign twiddle[86]  = 32'h3F176F5E; // cos: 0.492898, sin:0.870087
    assign twiddle[87]  = 32'h3DB87022; // cos: 0.482184, sin:0.876070
    assign twiddle[88]  = 32'h3C5670E2; // cos: 0.471397, sin:0.881921
    assign twiddle[89]  = 32'h3AF2719D; // cos: 0.460539, sin:0.887640
    assign twiddle[90]  = 32'h398C7254; // cos: 0.449611, sin:0.893224
    assign twiddle[91]  = 32'h38247307; // cos: 0.438616, sin:0.898674
    assign twiddle[92]  = 32'h36BA73B5; // cos: 0.427555, sin:0.903989
    assign twiddle[93]  = 32'h354D745F; // cos: 0.416430, sin:0.909168
    assign twiddle[94]  = 32'h33DF7504; // cos: 0.405241, sin:0.914210
    assign twiddle[95]  = 32'h326E75A5; // cos: 0.393992, sin:0.919114
    assign twiddle[96]  = 32'h30FB7641; // cos: 0.382683, sin:0.923880
    assign twiddle[97]  = 32'h2F8776D8; // cos: 0.371317, sin:0.928506
    assign twiddle[98]  = 32'h2E11776B; // cos: 0.359895, sin:0.932993
    assign twiddle[99]  = 32'h2C9977FA; // cos: 0.348419, sin:0.937339
    assign twiddle[100] = 32'h2B1F7884; // cos: 0.336890, sin:0.941544
    assign twiddle[101] = 32'h29A37909; // cos: 0.325310, sin:0.945607
    assign twiddle[102] = 32'h28267989; // cos: 0.313682, sin:0.949528
    assign twiddle[103] = 32'h26A87A05; // cos: 0.302006, sin:0.953306
    assign twiddle[104] = 32'h25287A7C; // cos: 0.290285, sin:0.956940
    assign twiddle[105] = 32'h23A67AEE; // cos: 0.278520, sin:0.960431
    assign twiddle[106] = 32'h22237B5C; // cos: 0.266713, sin:0.963776
    assign twiddle[107] = 32'h209F7BC5; // cos: 0.254866, sin:0.966976
    assign twiddle[108] = 32'h1F1A7C29; // cos: 0.242980, sin:0.970031
    assign twiddle[109] = 32'h1D937C88; // cos: 0.231058, sin:0.972940
    assign twiddle[110] = 32'h1C0B7CE3; // cos: 0.219101, sin:0.975702
    assign twiddle[111] = 32'h1A827D39; // cos: 0.207111, sin:0.978317
    assign twiddle[112] = 32'h18F97D89; // cos: 0.195090, sin:0.980785
    assign twiddle[113] = 32'h176E7DD5; // cos: 0.183040, sin:0.983105
    assign twiddle[114] = 32'h15E27E1D; // cos: 0.170962, sin:0.985278
    assign twiddle[115] = 32'h14557E5F; // cos: 0.158858, sin:0.987301
    assign twiddle[116] = 32'h12C87E9C; // cos: 0.146730, sin:0.989177
    assign twiddle[117] = 32'h113A7ED5; // cos: 0.134581, sin:0.990903
    assign twiddle[118] = 32'h0FAB7F09; // cos: 0.122411, sin:0.992480
    assign twiddle[119] = 32'h0E1C7F37; // cos: 0.110222, sin:0.993907
    assign twiddle[120] = 32'h0C8C7F61; // cos: 0.098017, sin:0.995185
    assign twiddle[121] = 32'h0AFB7F86; // cos: 0.085797, sin:0.996313
    assign twiddle[122] = 32'h096A7FA6; // cos: 0.073565, sin:0.997290
    assign twiddle[123] = 32'h07D97FC1; // cos: 0.061321, sin:0.998118
    assign twiddle[124] = 32'h06487FD8; // cos: 0.049068, sin:0.998795
    assign twiddle[125] = 32'h04B67FE9; // cos: 0.036807, sin:0.999322
    assign twiddle[126] = 32'h03247FF5; // cos: 0.024541, sin:0.999699
    assign twiddle[127] = 32'h01927FFD; // cos: 0.012272, sin:0.999925
    assign twiddle[128] = 32'h00007FFF; // cos: 0.000000, sin:1.000000
    assign twiddle[129] = 32'hFE6E7FFD; // cos: -0.012272, sin:0.999925
    assign twiddle[130] = 32'hFCDC7FF5; // cos: -0.024541, sin:0.999699
    assign twiddle[131] = 32'hFB4A7FE9; // cos: -0.036807, sin:0.999322
    assign twiddle[132] = 32'hF9B87FD8; // cos: -0.049068, sin:0.998795
    assign twiddle[133] = 32'hF8277FC1; // cos: -0.061321, sin:0.998118
    assign twiddle[134] = 32'hF6967FA6; // cos: -0.073565, sin:0.997290
    assign twiddle[135] = 32'hF5057F86; // cos: -0.085797, sin:0.996313
    assign twiddle[136] = 32'hF3747F61; // cos: -0.098017, sin:0.995185
    assign twiddle[137] = 32'hF1E47F37; // cos: -0.110222, sin:0.993907
    assign twiddle[138] = 32'hF0557F09; // cos: -0.122411, sin:0.992480
    assign twiddle[139] = 32'hEEC67ED5; // cos: -0.134581, sin:0.990903
    assign twiddle[140] = 32'hED387E9C; // cos: -0.146730, sin:0.989177
    assign twiddle[141] = 32'hEBAB7E5F; // cos: -0.158858, sin:0.987301
    assign twiddle[142] = 32'hEA1E7E1D; // cos: -0.170962, sin:0.985278
    assign twiddle[143] = 32'hE8927DD5; // cos: -0.183040, sin:0.983105
    assign twiddle[144] = 32'hE7077D89; // cos: -0.195090, sin:0.980785
    assign twiddle[145] = 32'hE57E7D39; // cos: -0.207111, sin:0.978317
    assign twiddle[146] = 32'hE3F57CE3; // cos: -0.219101, sin:0.975702
    assign twiddle[147] = 32'hE26D7C88; // cos: -0.231058, sin:0.972940
    assign twiddle[148] = 32'hE0E67C29; // cos: -0.242980, sin:0.970031
    assign twiddle[149] = 32'hDF617BC5; // cos: -0.254866, sin:0.966976
    assign twiddle[150] = 32'hDDDD7B5C; // cos: -0.266713, sin:0.963776
    assign twiddle[151] = 32'hDC5A7AEE; // cos: -0.278520, sin:0.960431
    assign twiddle[152] = 32'hDAD87A7C; // cos: -0.290285, sin:0.956940
    assign twiddle[153] = 32'hD9587A05; // cos: -0.302006, sin:0.953306
    assign twiddle[154] = 32'hD7DA7989; // cos: -0.313682, sin:0.949528
    assign twiddle[155] = 32'hD65D7909; // cos: -0.325310, sin:0.945607
    assign twiddle[156] = 32'hD4E17884; // cos: -0.336890, sin:0.941544
    assign twiddle[157] = 32'hD36777FA; // cos: -0.348419, sin:0.937339
    assign twiddle[158] = 32'hD1EF776B; // cos: -0.359895, sin:0.932993
    assign twiddle[159] = 32'hD07976D8; // cos: -0.371317, sin:0.928506
    assign twiddle[160] = 32'hCF057641; // cos: -0.382683, sin:0.923880
    assign twiddle[161] = 32'hCD9275A5; // cos: -0.393992, sin:0.919114
    assign twiddle[162] = 32'hCC217504; // cos: -0.405241, sin:0.914210
    assign twiddle[163] = 32'hCAB3745F; // cos: -0.416430, sin:0.909168
    assign twiddle[164] = 32'hC94673B5; // cos: -0.427555, sin:0.903989
    assign twiddle[165] = 32'hC7DC7307; // cos: -0.438616, sin:0.898674
    assign twiddle[166] = 32'hC6747254; // cos: -0.449611, sin:0.893224
    assign twiddle[167] = 32'hC50E719D; // cos: -0.460539, sin:0.887640
    assign twiddle[168] = 32'hC3AA70E2; // cos: -0.471397, sin:0.881921
    assign twiddle[169] = 32'hC2487022; // cos: -0.482184, sin:0.876070
    assign twiddle[170] = 32'hC0E96F5E; // cos: -0.492898, sin:0.870087
    assign twiddle[171] = 32'hBF8D6E96; // cos: -0.503538, sin:0.863973
    assign twiddle[172] = 32'hBE326DC9; // cos: -0.514103, sin:0.857729
    assign twiddle[173] = 32'hBCDB6CF8; // cos: -0.524590, sin:0.851355
    assign twiddle[174] = 32'hBB866C23; // cos: -0.534998, sin:0.844854
    assign twiddle[175] = 32'hBA336B4A; // cos: -0.545325, sin:0.838225
    assign twiddle[176] = 32'hB8E46A6D; // cos: -0.555570, sin:0.831470
    assign twiddle[177] = 32'hB797698B; // cos: -0.565732, sin:0.824589
    assign twiddle[178] = 32'hB64C68A6; // cos: -0.575808, sin:0.817585
    assign twiddle[179] = 32'hB50567BC; // cos: -0.585798, sin:0.810457
    assign twiddle[180] = 32'hB3C166CF; // cos: -0.595699, sin:0.803208
    assign twiddle[181] = 32'hB27F65DD; // cos: -0.605511, sin:0.795837
    assign twiddle[182] = 32'hB14164E8; // cos: -0.615232, sin:0.788346
    assign twiddle[183] = 32'hB00563EE; // cos: -0.624859, sin:0.780737
    assign twiddle[184] = 32'hAECD62F1; // cos: -0.634393, sin:0.773010
    assign twiddle[185] = 32'hAD9861F0; // cos: -0.643832, sin:0.765167
    assign twiddle[186] = 32'hAC6560EB; // cos: -0.653173, sin:0.757209
    assign twiddle[187] = 32'hAB375FE3; // cos: -0.662416, sin:0.749136
    assign twiddle[188] = 32'hAA0B5ED7; // cos: -0.671559, sin:0.740951
    assign twiddle[189] = 32'hA8E35DC7; // cos: -0.680601, sin:0.732654
    assign twiddle[190] = 32'hA7BE5CB3; // cos: -0.689541, sin:0.724247
    assign twiddle[191] = 32'hA69C5B9C; // cos: -0.698376, sin:0.715731
    assign twiddle[192] = 32'hA57E5A82; // cos: -0.707107, sin:0.707107
    assign twiddle[193] = 32'hA4645964; // cos: -0.715731, sin:0.698376
    assign twiddle[194] = 32'hA34D5842; // cos: -0.724247, sin:0.689541
    assign twiddle[195] = 32'hA239571D; // cos: -0.732654, sin:0.680601
    assign twiddle[196] = 32'hA12955F5; // cos: -0.740951, sin:0.671559
    assign twiddle[197] = 32'hA01D54C9; // cos: -0.749136, sin:0.662416
    assign twiddle[198] = 32'h9F15539B; // cos: -0.757209, sin:0.653173
    assign twiddle[199] = 32'h9E105268; // cos: -0.765167, sin:0.643832
    assign twiddle[200] = 32'h9D0F5133; // cos: -0.773010, sin:0.634393
    assign twiddle[201] = 32'h9C124FFB; // cos: -0.780737, sin:0.624859
    assign twiddle[202] = 32'h9B184EBF; // cos: -0.788346, sin:0.615232
    assign twiddle[203] = 32'h9A234D81; // cos: -0.795837, sin:0.605511
    assign twiddle[204] = 32'h99314C3F; // cos: -0.803208, sin:0.595699
    assign twiddle[205] = 32'h98444AFB; // cos: -0.810457, sin:0.585798
    assign twiddle[206] = 32'h975A49B4; // cos: -0.817585, sin:0.575808
    assign twiddle[207] = 32'h96754869; // cos: -0.824589, sin:0.565732
    assign twiddle[208] = 32'h9593471C; // cos: -0.831470, sin:0.555570
    assign twiddle[209] = 32'h94B645CD; // cos: -0.838225, sin:0.545325
    assign twiddle[210] = 32'h93DD447A; // cos: -0.844854, sin:0.534998
    assign twiddle[211] = 32'h93084325; // cos: -0.851355, sin:0.524590
    assign twiddle[212] = 32'h923741CE; // cos: -0.857729, sin:0.514103
    assign twiddle[213] = 32'h916A4073; // cos: -0.863973, sin:0.503538
    assign twiddle[214] = 32'h90A23F17; // cos: -0.870087, sin:0.492898
    assign twiddle[215] = 32'h8FDE3DB8; // cos: -0.876070, sin:0.482184
    assign twiddle[216] = 32'h8F1E3C56; // cos: -0.881921, sin:0.471397
    assign twiddle[217] = 32'h8E633AF2; // cos: -0.887640, sin:0.460539
    assign twiddle[218] = 32'h8DAC398C; // cos: -0.893224, sin:0.449611
    assign twiddle[219] = 32'h8CF93824; // cos: -0.898674, sin:0.438616
    assign twiddle[220] = 32'h8C4B36BA; // cos: -0.903989, sin:0.427555
    assign twiddle[221] = 32'h8BA1354D; // cos: -0.909168, sin:0.416430
    assign twiddle[222] = 32'h8AFC33DF; // cos: -0.914210, sin:0.405241
    assign twiddle[223] = 32'h8A5B326E; // cos: -0.919114, sin:0.393992
    assign twiddle[224] = 32'h89BF30FB; // cos: -0.923880, sin:0.382683
    assign twiddle[225] = 32'h89282F87; // cos: -0.928506, sin:0.371317
    assign twiddle[226] = 32'h88952E11; // cos: -0.932993, sin:0.359895
    assign twiddle[227] = 32'h88062C99; // cos: -0.937339, sin:0.348419
    assign twiddle[228] = 32'h877C2B1F; // cos: -0.941544, sin:0.336890
    assign twiddle[229] = 32'h86F729A3; // cos: -0.945607, sin:0.325310
    assign twiddle[230] = 32'h86772826; // cos: -0.949528, sin:0.313682
    assign twiddle[231] = 32'h85FB26A8; // cos: -0.953306, sin:0.302006
    assign twiddle[232] = 32'h85842528; // cos: -0.956940, sin:0.290285
    assign twiddle[233] = 32'h851223A6; // cos: -0.960431, sin:0.278520
    assign twiddle[234] = 32'h84A42223; // cos: -0.963776, sin:0.266713
    assign twiddle[235] = 32'h843B209F; // cos: -0.966976, sin:0.254866
    assign twiddle[236] = 32'h83D71F1A; // cos: -0.970031, sin:0.242980
    assign twiddle[237] = 32'h83781D93; // cos: -0.972940, sin:0.231058
    assign twiddle[238] = 32'h831D1C0B; // cos: -0.975702, sin:0.219101
    assign twiddle[239] = 32'h82C71A82; // cos: -0.978317, sin:0.207111
    assign twiddle[240] = 32'h827718F9; // cos: -0.980785, sin:0.195090
    assign twiddle[241] = 32'h822B176E; // cos: -0.983105, sin:0.183040
    assign twiddle[242] = 32'h81E315E2; // cos: -0.985278, sin:0.170962
    assign twiddle[243] = 32'h81A11455; // cos: -0.987301, sin:0.158858
    assign twiddle[244] = 32'h816412C8; // cos: -0.989177, sin:0.146730
    assign twiddle[245] = 32'h812B113A; // cos: -0.990903, sin:0.134581
    assign twiddle[246] = 32'h80F70FAB; // cos: -0.992480, sin:0.122411
    assign twiddle[247] = 32'h80C90E1C; // cos: -0.993907, sin:0.110222
    assign twiddle[248] = 32'h809F0C8C; // cos: -0.995185, sin:0.098017
    assign twiddle[249] = 32'h807A0AFB; // cos: -0.996313, sin:0.085797
    assign twiddle[250] = 32'h805A096A; // cos: -0.997290, sin:0.073565
    assign twiddle[251] = 32'h803F07D9; // cos: -0.998118, sin:0.061321
    assign twiddle[252] = 32'h80280648; // cos: -0.998795, sin:0.049068
    assign twiddle[253] = 32'h801704B6; // cos: -0.999322, sin:0.036807
    assign twiddle[254] = 32'h800B0324; // cos: -0.999699, sin:0.024541
    assign twiddle[255] = 32'h80030192; // cos: -0.999925, sin:0.012272

  assign twiddle_out = twiddle[twiddle_adr[7:0]];

endmodule
